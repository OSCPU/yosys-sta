// add the ram module for blackbox



